module TheLime();

endmodule