module Data(
    input wire [2:0] input_reg_readA_address, // 3-bit address for reading Operand A.
    input wire [2:0] input_reg_readB_address, // 3-bit address for reading Operand B.
	input wire input_reg_write, // Single-bit signal to enable write operation.
    input wire [15:0] input_reg_write_value, // 16-bit value for write operation.
    input wire [2:0] input_reg_write_address, // 3-bit address for write operation.
	input wire CLK, // Single-bit clock signal for synchronization.
    
    input wire [15:0] input_imm, // 16-bit input of the instruction for the immediate to be parsed
    input wire output_MDR, //mdr output
    
    output reg [15:0] output_imm // 16-bit output representing the immediate value generated by the Immediate Generator.
    output reg [15:0] output_reg_A, // 16-bit output representing data read from Register A.
    output reg [15:0] output_reg_B // 16-bit output representing data read from Register B.
  
);

    //mdr inst needs to come in

    ProgrammableRegisterFile register_inst (
    .clk(clk),
      .Output_IR_RegA(Output_IR_RegA),
      .Output_IR_RegB(Output_IR_RegB),
      .Output_IR_RegD(Output_IR_RegD),
      .Output_IR_Imm(Output_IR_Imm),
        .output_MDR(output_MDR),
            
    );


     
        
        
        .Output_memToReg(Output_memToReg),
      .output_reWrite(output_reWrite),
      .output_mem_data(output_mem_data),
      .output_ALU(output_ALU),
      .input_imm(input_imm),
      
      .output_imm(output_imm),
      .output_reg_A(output_reg_A),
      .output_reg_B(output_reg_B),
      

    
endmodule
