
/*
 Author: Tulsi Manohar
 Date: 2/7/2024

 edited: 2/15/2024
*/

module Data(
    input wire [2:0] input_reg_readA_address, // 3-bit address for reading Operand A.
    input wire [2:0] input_reg_readB_address, // 3-bit address for reading Operand B.
    input wire input_reg_write, // Single-bit signal to enable write operation.
    input wire [2:0] input_reg_write_address, // 3-bit address for write operation.
    input wire CLK, // Single-bit clock signal for synchronization.
    input wire [15:0] input_imm, // 16-bit input of the instruction for the immediate to be parsed
    input wire input_branch,
    input wire [15:0] input_ALUOut,
    input wire [15:0] input_MDR,
    input wire memToReg,
    output wire [15:0] output_imm, // 16-bit output representing the immediate value generated by the Immediate Generator.
    output wire [15:0] output_reg_A, // 16-bit output representing data read from Register A.
    output wire [15:0] output_reg_B // 16-bit output representing data read from Register B.
);

reg [15:0] BorRd;
always @(*) begin
    case(input_branch)
        0: BorRd = input_reg_readB_address;
        1: BorRd = input_reg_write_address; 
        default: BorRd = 16'b0000_0000_0000_0000; // Default to zero if an invalid selection
    endcase
end

wire[15:0] registerInput;
mux2to1 IorD(
	.a(input_ALUOut),
	.b(input_MDR),
	.select(memToReg),
	.out(registerInput)
);

ProgrammableRegisterFile register_inst (
    .CLK(CLK),
    .input_reg_readA_address(input_reg_readA_address),
    .input_reg_readB_address(BorRd),
    .input_reg_write(input_reg_write),
    .input_reg_write_value(registerInput), // Changed from 'immOrOut'
    .input_reg_write_address(input_reg_write_address),
    .output_reg_A(output_reg_A),
    .output_reg_B(output_reg_B)
);

ImmediateGenerator ig_inst(
    .input_imm(input_imm),
    .output_imm(output_imm)
);



endmodule
