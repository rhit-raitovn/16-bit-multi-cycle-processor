module Data(
    input wire clk,
    input wire [6:0] Output_IR_Control, // 7-bit output for opcode and func4.
    input wire [3:0] Output_IR_RegA, // 3-bit output for register A address.
    input wire [3:0] Output_IR_RegB, // 3-bit output for register B address.
    input wire [3:0] Output_IR_RegD, // 3-bit output for register D address.
    input wire [15:0] Output_IR_Imm, // 16-bit output for immediate value.
    input wire [0:0] Output_memToReg, output_regWrite,
    input wire [15:0] output_MDR,
    input wire [15:0] output_ALU,
    input wire [15:0] input_imm, // 16-bit input of the instruction for the immediate to be parsed


  
    output reg [15:0] output_imm, // 16-bit output representing the immediate value generated by the Immediate Generator.
    output reg [15:0] output_reg_A, // 16-bit output representing data read from Register A.
    output reg [15:0] output_reg_B // 16-bit output representing data read from Register B.
  
);

    //mdr inst needs to come in

    ProgrammableRegisterFile register_inst (
    .clk(clk),
      .Output_IR_RegA(Output_IR_RegA),
      .Output_IR_RegB(Output_IR_RegB),
      .Output_IR_RegD(Output_IR_RegD),
      .Output_IR_Imm(Output_IR_Imm),
        .output_MDR(output_MDR),
            
    );


     
        
        
        .Output_memToReg(Output_memToReg),
      .output_reWrite(output_reWrite),
      .output_mem_data(output_mem_data),
      .output_ALU(output_ALU),
      .input_imm(input_imm),
      
      .output_imm(output_imm),
      .output_reg_A(output_reg_A),
      .output_reg_B(output_reg_B),
      

    
endmodule
