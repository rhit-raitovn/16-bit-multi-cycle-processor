module Data(
    	input wire [2:0] input_reg_readA_address, // 3-bit address for reading Operand A.
    	input wire [2:0] input_reg_readB_address, // 3-bit address for reading Operand B.
	input wire input_reg_write, // Single-bit signal to enable write operation.
    	input wire [2:0] input_reg_write_address, // 3-bit address for write operation.
	input wire CLK, // Single-bit clock signal for synchronization.
    
    	input wire [15:0] input_imm, // 16-bit input of the instruction for the immediate to be parsed

	input wire [15:0] input_ALUOut,
	input wire [15:0] input_MDR,
  	input wire memToReg,
  
	
	output wire [15:0] output_imm, // 16-bit output representing the immediate value generated by the Immediate Generator.
    output wire [15:0] output_reg_A, // 16-bit output representing data read from Register A.
    output wire [15:0] output_reg_B // 16-bit output representing data read from Register B.
  
);


    ProgrammableRegisterFile register_inst (
	    
	    .CLK(CLK),
	    .input_reg_readA_address(input_reg_readA_address),
	    .input_reg_readB_address(input_reg_readB_address),
	    .input_reg_write(input_reg_write),
	    .input_reg_write_value(immOrOut),
	    .input_reg_write_address(input_reg_write_address),
	    .output_reg_A(output_reg_A),
	    .output_reg_B(output_reg_B)
   	);

	ImmediateGenerator ig_inst(
	    .input_imm(input_imm),
	    .output_imm(output_imm)
	);
         
	
	reg [15:0] immOrOut;
	mux2to1 mux_inst(
		.a(input_ALUOut),
		.b(input_MDR),
		.select(memToReg),
		.out(immOrOut)
	);

    
endmodule
